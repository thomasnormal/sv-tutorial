module adder(
  input  logic [7:0] a,
  input  logic [7:0] b,
  output logic [7:0] sum
);
  // TODO: drive sum combinationally from a and b
endmodule
