module adder (
  input  logic [3:0] A, B,
  output logic [4:0] X
);
  // TODO: compute X as the sum of A and B
endmodule
