module top;
  initial begin
    // TODO: print a greeting with $display, then call $finish
  end
endmodule
