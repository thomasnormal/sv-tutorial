module top;
  initial begin
    $display("Hello, SRAM world!");
    $finish;
  end
endmodule
