interface adder_if (input logic clk);
  logic [7:0] a, b, sum;
  logic       carry;
endinterface
