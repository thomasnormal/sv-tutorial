module top;
  initial begin
    // TODO: $display("hello, world");
  end
endmodule
