// A packed struct maps named fields onto a contiguous bit-vector.
// Fields are declared MSB-first; we need we, addr, and wdata.
package mem_pkg;
  typedef struct packed {
    // TODO: add the three fields of the SRAM command bus
  } mem_cmd_t;
endpackage
